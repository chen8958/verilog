module tb ();

initial begin
  $display("hello vcs");
end

endmodule